`default_nettype none

//`define NO_MUACM
//`define SPI_DRIVEN
`define BUS_DRIVEN

module sid_clk(
    input CLK,
    output CLKen
    );

  reg [4:0] counter;
  wire CLKen = (counter == 0);

  initial begin
      counter <= 0;
  end

  always @(posedge CLK) begin
      if (CLKen) begin
          counter <= 5'd23;
      end else begin
          counter <= counter - 5'd1;
      end
  end
endmodule

// A very crappy filter
// y(n) = y(n-1) * 7/8 + x(n)
module simple_filter(
    input                CLK,
    input                CLKen,
    input  signed [15:0] in,
    output signed [15:0] out,
    );

  reg signed [21:0] accum;
  assign out = accum[20:5];

  initial begin
    accum <= 0;
  end

  always @(posedge CLK) begin
    if (CLKen) begin
      accum <= (accum - (accum >>> 3)) + in;
    end
  end
endmodule

module top (
    // I2S
    output wire i2s_din,
    input  wire i2s_dout,
    input  wire i2s_sclk,
    input  wire i2s_lrclk,
    // I2C (shared)
    inout  wire scl_led,
    inout  wire sda_btn,
    // USB
    inout  wire usb_dp,
    inout  wire usb_dn,
    output wire usb_pu,
    // Clock
    input  wire sys_clk,
`ifdef SPI_DRIVEN
    // SPI bus
    input wire d0,  // SCLK
    input wire d1,  // MOSI
    input wire d2   // CS
`endif
`ifdef BUS_DRIVEN
    // data bus
    inout  wire d0,
    inout  wire d1,
    inout  wire d2,
    inout  wire d3,
    inout  wire d4,
    inout  wire d5,
    inout  wire d6,
    inout  wire d7,
    // address bus
    inout  wire a0,
    inout  wire a1,
    inout  wire a2,
    inout  wire a3,
    inout  wire a4,
    // sid clock
    inout  wire phi2,
    // sid chip select
    inout  wire cs_n,
    // sid read/write
    inout  wire rw
`endif
);

`ifdef SPI_DRIVEN
    // SPI slave
    reg [7:0] spi_data;
    reg spi_recv;
    spi_slave spi(
        sys_clk,            // system clock
        d0,                 // spi clock
        d1,                 // spi mosi
        d2,                 // spi chip select
        spi_data,           // data out
        spi_recv            // data received
    );

    // input data decoder
    //
    // receive format:
    //    1AAA AADD   - address, data MSB
    //    0?DD DDDD   -          data LSB
    //
    reg [4:0] addrBusIn;    // latched address
    reg [7:0] dataBusIn;    // latched data
    reg wrStrobe;           // write signal
    always @(posedge sys_clk) begin
        if (spi_recv) begin
            if (spi_data[7] == 'b1) begin
                wrStrobe <= 0;
                addrBusIn <= spi_data[6:2];
                dataBusIn <= { spi_data[1:0], dataBusIn[5:0] };
            end else begin
                wrStrobe <= 1;
                dataBusIn <= { dataBusIn[7:6], spi_data[5:0] };
            end
        end else begin
            wrStrobe <= 0;
        end
    end

    // SID 1Mhz clock
    wire CLKen;
    sid_clk sid_clk_en(sys_clk, CLKen);
`endif
`ifdef BUS_DRIVEN

    reg        wrStrobe;
    reg        dataBusOE;
    reg  [7:0] dataBusOut;
    wire [7:0] dataBusIn;
    wire [4:0] addrBusIn;

    wire sidCLK, sidCS, sidRW;

    initial begin
        dataBusOE  <= 0;
        dataBusOut <= 0;
        sidCLKPrev <= 0;
        wrStrobe   <= 0;
    end

    SB_IO #(
        .PIN_TYPE(6'b1010_00),  // Reg input, tristate output
        .PULLUP(1'b0)
    ) dataBusPins[7:0] (
        .PACKAGE_PIN({d7, d6, d5, d4, d3, d2, d1, d0}),
        .OUTPUT_ENABLE({8{ dataBusOE }}),
        .INPUT_CLK(sys_clk),
        .D_OUT_0(dataBusOut),
        .D_IN_0(dataBusIn)
    );

    SB_IO #(
        .PIN_TYPE(6'b0000_00),  // Reg input, no output
        .PULLUP(1'b0),
    ) addrBusPins[4:0] (
        .PACKAGE_PIN({a4, a3, a2, a1, a0}),
        .INPUT_CLK(sys_clk),
        .D_IN_0(addrBusIn)
    );

    SB_IO #(
        .PIN_TYPE(6'b0000_00),  // Reg input, no output
        .PULLUP(1'b0)
    ) ctrlBusPins[2:0] (
        .PACKAGE_PIN({ phi2, cs_n, rw }),
        .INPUT_CLK(sys_clk),
        .D_IN_0({sidCLK, sidCS, sidRW})
    );

    reg CLKen;
    reg sidCLKPrev;
    always @(posedge sys_clk) begin
        sidCLKPrev <= sidCLK;
        CLKen      <= (sidCLKPrev & !sidCLK);
        wrStrobe   <= (sidCLKPrev & !sidCLK) & !sidCS & !sidRW;
    end
`endif

    wire signed [15:0] flt_out;
    simple_filter flt(sys_clk, CLKen, sid_out, flt_out);

    // SID
    wire signed [15:0] sid_out;
    sid the_sid(
           sys_clk,             // Master clock
           CLKen,               // 1Mhz enable
           wrStrobe,            // write data to sid addr
           addrBusIn,
           dataBusIn,
           sid_out);

    // I2S encoder
    wire i2s_sampled;
    i2s i2s_tx(
        sys_clk,
        flt_out,
        i2s_sclk,
        i2s_lrclk,
        i2s_din,
        i2s_sampled
    );

    // Little blinky
    wire led = CLKen;

    // I2C setup
    i2c_state_machine ism(
        .scl_led(scl_led),
        .sda_btn(sda_btn),
        .btn    (),
        .led    (led),
        .done   (),
        .clk    (sys_clk),
        .rst    (rst)
    );

`ifndef NO_MUACM
    // Local signals
    wire bootloader;
    reg boot = 1'b0;

    // Instance
    muacm acm_I(
        .usb_dp       (usb_dp),
        .usb_dn       (usb_dn),
        .usb_pu       (usb_pu),
        .in_data      (8'h00),
        .in_last      (),
        .in_valid     (1'b0),
        .in_ready     (),
        .in_flush_now (1'b0),
        .in_flush_time(1'b1),
        .out_data     (),
        .out_last     (),
        .out_valid    (),
        .out_ready    (1'b1),
        .bootloader   (bootloader),
        .clk          (clk_usb),
        .rst          (rst_usb)
    );

    // Warmboot
    always @(posedge clk_usb) begin
        boot <= boot | bootloader;
    end

    SB_WARMBOOT warmboot(
        .BOOT (boot),
        .S0   (1'b1),
        .S1   (1'b0)
    );
`endif

    // Local reset
    reg [15:0] rst_cnt = 0;
    wire rst_i = ~rst_cnt[15];
    always @(posedge sys_clk) begin
        if (~rst_cnt[15]) begin
            rst_cnt <= rst_cnt + 1;
        end
    end

    // Promote reset signal to global buffer
    wire rst;
    SB_GB rst_gbuf_I(
        .USER_SIGNAL_TO_GLOBAL_BUFFER(rst_i),
        .GLOBAL_BUFFER_OUTPUT(rst)
    );

    // Use HF OSC to generate USB clock
    wire clk_usb;
    wire rst_usb;
    sysmgr_hfosc sysmgr_I(
        .rst_in (rst),
        .clk_out(clk_usb),
        .rst_out(rst_usb)
    );
endmodule
